package shared_pkg;
    
    // Declare variables with data types
    integer test_finished=0;
    integer error_count=0;
    integer correct_count=0;

    function set_test_finish ();
        test_finished=1;
    endfunction

endpackage
